
import "DPI-C" function void info_reg(input logic[31:0] rf_data[] );
module RegisterFile #(ADDR_WIDTH = 5, DATA_WIDTH = 32) (
  input wire clk,
	input wire info_r,
  //写端口
  input wire wen,
  input wire [ADDR_WIDTH-1:0] waddr,
  input wire [DATA_WIDTH-1:0] wdata,
  //读端口1
  input  wire[ADDR_WIDTH-1:0] raddr1,
  output wire[DATA_WIDTH-1:0] rdata1
  //读端口2
  // input  wire[ADDR_WIDTH-1:0] raddr2,
  // output wire[DATA_WIDTH-1:0] rdata2
);

//寄存器
  reg [DATA_WIDTH-1:0] rf [2**ADDR_WIDTH-1:0];

//传出reg的值
always @(*)begin
	if(info_r == 1)begin
		info_reg(rf);
	end
end


//READ 1
assign rdata1 = (raddr1 == 5'b0) ? 32'b0 : rf[raddr1];

//READ 2
// assign rdata2 = (raddr2 == 5'b0) ? 32'b0 : rf[raddr2];

//WRITE
  always @(posedge clk) begin
    if(wen && waddr!=5'b0) rf[waddr] <= wdata;
  end



endmodule

